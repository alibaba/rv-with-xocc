/* 
*Copyright (c) 2021, Alibaba Group;
*Licensed under the Apache License, Version 2.0 (the "License");
*you may not use this file except in compliance with the License.
*You may obtain a copy of the License at

*   http://www.apache.org/licenses/LICENSE-2.0

*Unless required by applicable law or agreed to in writing, software
*distributed under the License is distributed on an "AS IS" BASIS,
*WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
*See the License for the specific language governing permissions and
*limitations under the License.
*/

// &ModuleBeg; @1
module soc_top(
  rv_0_clk,
  rv_0_retire_pc,
  rv_0_rst_addr,
  rv_0_rstn,
  dsa_0_clk,
  dsa_0_rstn,
  dsa_1_clk,
  dsa_1_rstn,
  dsa_2_clk,
  dsa_2_rstn,
  mem_sub_sys_clk,
  mem_sub_sys_rstn,
  rv_1_clk,
  rv_1_retire_pc,
  rv_1_rst_addr,
  rv_1_rstn,
  rv_2_clk,
  rv_2_retire_pc,
  rv_2_rst_addr,
  rv_2_rstn
);

// &Ports; @2
input             rv_0_clk;              
input   [31  :0]  rv_0_rst_addr;         
input             rv_0_rstn;             
input             dsa_0_clk;                   
input             dsa_0_rstn;                  
input             dsa_1_clk;                   
input             dsa_1_rstn;                  
input             dsa_2_clk;                   
input             dsa_2_rstn;                  
input             mem_sub_sys_clk;             
input             mem_sub_sys_rstn;            
input             rv_1_clk;               
input   [31  :0]  rv_1_rst_addr;          
input             rv_1_rstn;              
input             rv_2_clk;               
input   [31  :0]  rv_2_rst_addr;          
input             rv_2_rstn;              
output  [31  :0]  rv_0_retire_pc;        
output  [31  :0]  rv_1_retire_pc;         
output  [31  :0]  rv_2_retire_pc;         

// &Regs; @3

// &Wires; @4
wire              rv_0_clk;              
wire    [31  :0]  rv_0_m_axi_araddr;     
wire    [1   :0]  rv_0_m_axi_arburst;    
wire    [3   :0]  rv_0_m_axi_arcache;    
wire    [3   :0]  rv_0_m_axi_arid;       
wire    [7   :0]  rv_0_m_axi_arlen;      
wire    [0   :0]  rv_0_m_axi_arlock;     
wire    [2   :0]  rv_0_m_axi_arprot;     
wire    [3   :0]  rv_0_m_axi_arqos;      
wire              rv_0_m_axi_arready;    
wire    [2   :0]  rv_0_m_axi_arsize;     
wire              rv_0_m_axi_arvalid;    
wire    [31  :0]  rv_0_m_axi_awaddr;     
wire    [1   :0]  rv_0_m_axi_awburst;    
wire    [3   :0]  rv_0_m_axi_awcache;    
wire    [3   :0]  rv_0_m_axi_awid;       
wire    [7   :0]  rv_0_m_axi_awlen;      
wire    [0   :0]  rv_0_m_axi_awlock;     
wire    [2   :0]  rv_0_m_axi_awprot;     
wire    [3   :0]  rv_0_m_axi_awqos;      
wire              rv_0_m_axi_awready;    
wire    [2   :0]  rv_0_m_axi_awsize;     
wire              rv_0_m_axi_awvalid;    
wire    [3   :0]  rv_0_m_axi_bid;        
wire              rv_0_m_axi_bready;     
wire    [1   :0]  rv_0_m_axi_bresp;      
wire              rv_0_m_axi_bvalid;     
wire    [31  :0]  rv_0_m_axi_rdata;      
wire    [3   :0]  rv_0_m_axi_rid;        
wire              rv_0_m_axi_rlast;      
wire              rv_0_m_axi_rready;     
wire    [1   :0]  rv_0_m_axi_rresp;      
wire              rv_0_m_axi_rvalid;     
wire    [31  :0]  rv_0_m_axi_wdata;      
wire              rv_0_m_axi_wlast;      
wire              rv_0_m_axi_wready;     
wire    [3   :0]  rv_0_m_axi_wstrb;      
wire              rv_0_m_axi_wvalid;     
wire    [31  :0]  rv_0_retire_pc;        
wire    [31  :0]  rv_0_rst_addr;         
wire              rv_0_rstn;             
wire    [95  :0]  rv_0_xocc_2_cmd_buffer; 
wire              rv_0_xocc_2_cmd_empty; 
wire              rv_0_xocc_2_cmd_rd_en; 
wire    [31  :0]  rv_0_xocc_2_rsp_buffer; 
wire              rv_0_xocc_2_rsp_full;  
wire              rv_0_xocc_2_rsp_wr_en; 
wire              dsa_0_clk;                   
wire    [31  :0]  dsa_0_m_axi_araddr;          
wire    [1   :0]  dsa_0_m_axi_arburst;         
wire    [3   :0]  dsa_0_m_axi_arcache;         
wire    [3   :0]  dsa_0_m_axi_arid;            
wire    [7   :0]  dsa_0_m_axi_arlen;           
wire    [0   :0]  dsa_0_m_axi_arlock;          
wire    [2   :0]  dsa_0_m_axi_arprot;          
wire    [3   :0]  dsa_0_m_axi_arqos;           
wire              dsa_0_m_axi_arready;         
wire    [2   :0]  dsa_0_m_axi_arsize;          
wire              dsa_0_m_axi_arvalid;         
wire    [31  :0]  dsa_0_m_axi_awaddr;          
wire    [1   :0]  dsa_0_m_axi_awburst;         
wire    [3   :0]  dsa_0_m_axi_awcache;         
wire    [3   :0]  dsa_0_m_axi_awid;            
wire    [7   :0]  dsa_0_m_axi_awlen;           
wire    [0   :0]  dsa_0_m_axi_awlock;          
wire    [2   :0]  dsa_0_m_axi_awprot;          
wire    [3   :0]  dsa_0_m_axi_awqos;           
wire              dsa_0_m_axi_awready;         
wire    [2   :0]  dsa_0_m_axi_awsize;          
wire              dsa_0_m_axi_awvalid;         
wire    [3   :0]  dsa_0_m_axi_bid;             
wire              dsa_0_m_axi_bready;          
wire    [1   :0]  dsa_0_m_axi_bresp;           
wire              dsa_0_m_axi_bvalid;          
wire    [1023:0]  dsa_0_m_axi_rdata;           
wire    [3   :0]  dsa_0_m_axi_rid;             
wire              dsa_0_m_axi_rlast;           
wire              dsa_0_m_axi_rready;          
wire    [1   :0]  dsa_0_m_axi_rresp;           
wire              dsa_0_m_axi_rvalid;          
wire    [1023:0]  dsa_0_m_axi_wdata;           
wire              dsa_0_m_axi_wlast;           
wire              dsa_0_m_axi_wready;          
wire    [127 :0]  dsa_0_m_axi_wstrb;           
wire              dsa_0_m_axi_wvalid;          
wire              dsa_0_rstn;                  
wire              dsa_1_clk;                   
wire    [31  :0]  dsa_1_m_axi_araddr;          
wire    [1   :0]  dsa_1_m_axi_arburst;         
wire    [3   :0]  dsa_1_m_axi_arcache;         
wire    [3   :0]  dsa_1_m_axi_arid;            
wire    [7   :0]  dsa_1_m_axi_arlen;           
wire    [0   :0]  dsa_1_m_axi_arlock;          
wire    [2   :0]  dsa_1_m_axi_arprot;          
wire    [3   :0]  dsa_1_m_axi_arqos;           
wire              dsa_1_m_axi_arready;         
wire    [2   :0]  dsa_1_m_axi_arsize;          
wire              dsa_1_m_axi_arvalid;         
wire    [31  :0]  dsa_1_m_axi_awaddr;          
wire    [1   :0]  dsa_1_m_axi_awburst;         
wire    [3   :0]  dsa_1_m_axi_awcache;         
wire    [3   :0]  dsa_1_m_axi_awid;            
wire    [7   :0]  dsa_1_m_axi_awlen;           
wire    [0   :0]  dsa_1_m_axi_awlock;          
wire    [2   :0]  dsa_1_m_axi_awprot;          
wire    [3   :0]  dsa_1_m_axi_awqos;           
wire              dsa_1_m_axi_awready;         
wire    [2   :0]  dsa_1_m_axi_awsize;          
wire              dsa_1_m_axi_awvalid;         
wire    [3   :0]  dsa_1_m_axi_bid;             
wire              dsa_1_m_axi_bready;          
wire    [1   :0]  dsa_1_m_axi_bresp;           
wire              dsa_1_m_axi_bvalid;          
wire    [1023:0]  dsa_1_m_axi_rdata;           
wire    [3   :0]  dsa_1_m_axi_rid;             
wire              dsa_1_m_axi_rlast;           
wire              dsa_1_m_axi_rready;          
wire    [1   :0]  dsa_1_m_axi_rresp;           
wire              dsa_1_m_axi_rvalid;          
wire    [1023:0]  dsa_1_m_axi_wdata;           
wire              dsa_1_m_axi_wlast;           
wire              dsa_1_m_axi_wready;          
wire    [127 :0]  dsa_1_m_axi_wstrb;           
wire              dsa_1_m_axi_wvalid;          
wire              dsa_1_rstn;                  
wire              dsa_2_clk;                   
wire    [31  :0]  dsa_2_m_axi_araddr;          
wire    [1   :0]  dsa_2_m_axi_arburst;         
wire    [3   :0]  dsa_2_m_axi_arcache;         
wire    [3   :0]  dsa_2_m_axi_arid;            
wire    [7   :0]  dsa_2_m_axi_arlen;           
wire    [0   :0]  dsa_2_m_axi_arlock;          
wire    [2   :0]  dsa_2_m_axi_arprot;          
wire    [3   :0]  dsa_2_m_axi_arqos;           
wire              dsa_2_m_axi_arready;         
wire    [2   :0]  dsa_2_m_axi_arsize;          
wire              dsa_2_m_axi_arvalid;         
wire    [31  :0]  dsa_2_m_axi_awaddr;          
wire    [1   :0]  dsa_2_m_axi_awburst;         
wire    [3   :0]  dsa_2_m_axi_awcache;         
wire    [3   :0]  dsa_2_m_axi_awid;            
wire    [7   :0]  dsa_2_m_axi_awlen;           
wire    [0   :0]  dsa_2_m_axi_awlock;          
wire    [2   :0]  dsa_2_m_axi_awprot;          
wire    [3   :0]  dsa_2_m_axi_awqos;           
wire              dsa_2_m_axi_awready;         
wire    [2   :0]  dsa_2_m_axi_awsize;          
wire              dsa_2_m_axi_awvalid;         
wire    [3   :0]  dsa_2_m_axi_bid;             
wire              dsa_2_m_axi_bready;          
wire    [1   :0]  dsa_2_m_axi_bresp;           
wire              dsa_2_m_axi_bvalid;          
wire    [1023:0]  dsa_2_m_axi_rdata;           
wire    [3   :0]  dsa_2_m_axi_rid;             
wire              dsa_2_m_axi_rlast;           
wire              dsa_2_m_axi_rready;          
wire    [1   :0]  dsa_2_m_axi_rresp;           
wire              dsa_2_m_axi_rvalid;          
wire    [1023:0]  dsa_2_m_axi_wdata;           
wire              dsa_2_m_axi_wlast;           
wire              dsa_2_m_axi_wready;          
wire    [127 :0]  dsa_2_m_axi_wstrb;           
wire              dsa_2_m_axi_wvalid;          
wire              dsa_2_rstn;                  
wire              mem_sub_sys_clk;             
wire              mem_sub_sys_rstn;            
wire              rv_1_clk;               
wire    [31  :0]  rv_1_m_axi_araddr;      
wire    [1   :0]  rv_1_m_axi_arburst;     
wire    [3   :0]  rv_1_m_axi_arcache;     
wire    [3   :0]  rv_1_m_axi_arid;        
wire    [7   :0]  rv_1_m_axi_arlen;       
wire    [0   :0]  rv_1_m_axi_arlock;      
wire    [2   :0]  rv_1_m_axi_arprot;      
wire    [3   :0]  rv_1_m_axi_arqos;       
wire              rv_1_m_axi_arready;     
wire    [2   :0]  rv_1_m_axi_arsize;      
wire              rv_1_m_axi_arvalid;     
wire    [31  :0]  rv_1_m_axi_awaddr;      
wire    [1   :0]  rv_1_m_axi_awburst;     
wire    [3   :0]  rv_1_m_axi_awcache;     
wire    [3   :0]  rv_1_m_axi_awid;        
wire    [7   :0]  rv_1_m_axi_awlen;       
wire    [0   :0]  rv_1_m_axi_awlock;      
wire    [2   :0]  rv_1_m_axi_awprot;      
wire    [3   :0]  rv_1_m_axi_awqos;       
wire              rv_1_m_axi_awready;     
wire    [2   :0]  rv_1_m_axi_awsize;      
wire              rv_1_m_axi_awvalid;     
wire    [3   :0]  rv_1_m_axi_bid;         
wire              rv_1_m_axi_bready;      
wire    [1   :0]  rv_1_m_axi_bresp;       
wire              rv_1_m_axi_bvalid;      
wire    [31  :0]  rv_1_m_axi_rdata;       
wire    [3   :0]  rv_1_m_axi_rid;         
wire              rv_1_m_axi_rlast;       
wire              rv_1_m_axi_rready;      
wire    [1   :0]  rv_1_m_axi_rresp;       
wire              rv_1_m_axi_rvalid;      
wire    [31  :0]  rv_1_m_axi_wdata;       
wire              rv_1_m_axi_wlast;       
wire              rv_1_m_axi_wready;      
wire    [3   :0]  rv_1_m_axi_wstrb;       
wire              rv_1_m_axi_wvalid;      
wire    [31  :0]  rv_1_retire_pc;         
wire    [31  :0]  rv_1_rst_addr;          
wire              rv_1_rstn;              
wire    [95  :0]  rv_1_xocc_3_cmd_buffer; 
wire              rv_1_xocc_3_cmd_empty;  
wire              rv_1_xocc_3_cmd_rd_en;  
wire    [31  :0]  rv_1_xocc_3_rsp_buffer; 
wire              rv_1_xocc_3_rsp_full;   
wire              rv_1_xocc_3_rsp_wr_en;  
wire              rv_2_clk;               
wire    [31  :0]  rv_2_m_axi_araddr;      
wire    [1   :0]  rv_2_m_axi_arburst;     
wire    [3   :0]  rv_2_m_axi_arcache;     
wire    [3   :0]  rv_2_m_axi_arid;        
wire    [7   :0]  rv_2_m_axi_arlen;       
wire    [0   :0]  rv_2_m_axi_arlock;      
wire    [2   :0]  rv_2_m_axi_arprot;      
wire    [3   :0]  rv_2_m_axi_arqos;       
wire              rv_2_m_axi_arready;     
wire    [2   :0]  rv_2_m_axi_arsize;      
wire              rv_2_m_axi_arvalid;     
wire    [31  :0]  rv_2_m_axi_awaddr;      
wire    [1   :0]  rv_2_m_axi_awburst;     
wire    [3   :0]  rv_2_m_axi_awcache;     
wire    [3   :0]  rv_2_m_axi_awid;        
wire    [7   :0]  rv_2_m_axi_awlen;       
wire    [0   :0]  rv_2_m_axi_awlock;      
wire    [2   :0]  rv_2_m_axi_awprot;      
wire    [3   :0]  rv_2_m_axi_awqos;       
wire              rv_2_m_axi_awready;     
wire    [2   :0]  rv_2_m_axi_awsize;      
wire              rv_2_m_axi_awvalid;     
wire    [3   :0]  rv_2_m_axi_bid;         
wire              rv_2_m_axi_bready;      
wire    [1   :0]  rv_2_m_axi_bresp;       
wire              rv_2_m_axi_bvalid;      
wire    [31  :0]  rv_2_m_axi_rdata;       
wire    [3   :0]  rv_2_m_axi_rid;         
wire              rv_2_m_axi_rlast;       
wire              rv_2_m_axi_rready;      
wire    [1   :0]  rv_2_m_axi_rresp;       
wire              rv_2_m_axi_rvalid;      
wire    [31  :0]  rv_2_m_axi_wdata;       
wire              rv_2_m_axi_wlast;       
wire              rv_2_m_axi_wready;      
wire    [3   :0]  rv_2_m_axi_wstrb;       
wire              rv_2_m_axi_wvalid;      
wire    [31  :0]  rv_2_retire_pc;         
wire    [31  :0]  rv_2_rst_addr;          
wire              rv_2_rstn;              
wire    [95  :0]  rv_2_xocc_4_cmd_buffer; 
wire              rv_2_xocc_4_cmd_empty;  
wire              rv_2_xocc_4_cmd_rd_en;  
wire    [31  :0]  rv_2_xocc_4_rsp_buffer; 
wire              rv_2_xocc_4_rsp_full;   
wire              rv_2_xocc_4_rsp_wr_en;  
wire    [31  :0]  s_0_axi_araddr;              
wire    [1   :0]  s_0_axi_arburst;             
wire    [3   :0]  s_0_axi_arcache;             
wire    [7   :0]  s_0_axi_arid;                
wire    [7   :0]  s_0_axi_arlen;               
wire    [0   :0]  s_0_axi_arlock;              
wire    [2   :0]  s_0_axi_arprot;              
wire    [3   :0]  s_0_axi_arqos;               
wire              s_0_axi_arready;             
wire    [2   :0]  s_0_axi_arsize;              
wire              s_0_axi_arvalid;             
wire    [31  :0]  s_0_axi_awaddr;              
wire    [1   :0]  s_0_axi_awburst;             
wire    [3   :0]  s_0_axi_awcache;             
wire    [7   :0]  s_0_axi_awid;                
wire    [7   :0]  s_0_axi_awlen;               
wire    [0   :0]  s_0_axi_awlock;              
wire    [2   :0]  s_0_axi_awprot;              
wire    [3   :0]  s_0_axi_awqos;               
wire              s_0_axi_awready;             
wire    [2   :0]  s_0_axi_awsize;              
wire              s_0_axi_awvalid;             
wire    [7   :0]  s_0_axi_bid;                 
wire              s_0_axi_bready;              
wire    [1   :0]  s_0_axi_bresp;               
wire              s_0_axi_bvalid;              
wire    [1023:0]  s_0_axi_rdata;               
wire    [7   :0]  s_0_axi_rid;                 
wire              s_0_axi_rlast;               
wire              s_0_axi_rready;              
wire    [1   :0]  s_0_axi_rresp;               
wire              s_0_axi_rvalid;              
wire    [1023:0]  s_0_axi_wdata;               
wire              s_0_axi_wlast;               
wire              s_0_axi_wready;              
wire    [127 :0]  s_0_axi_wstrb;               
wire              s_0_axi_wvalid;              
wire    [31  :0]  s_1_axi_araddr;              
wire    [1   :0]  s_1_axi_arburst;             
wire    [3   :0]  s_1_axi_arcache;             
wire    [7   :0]  s_1_axi_arid;                
wire    [7   :0]  s_1_axi_arlen;               
wire    [0   :0]  s_1_axi_arlock;              
wire    [2   :0]  s_1_axi_arprot;              
wire    [3   :0]  s_1_axi_arqos;               
wire              s_1_axi_arready;             
wire    [2   :0]  s_1_axi_arsize;              
wire              s_1_axi_arvalid;             
wire    [31  :0]  s_1_axi_awaddr;              
wire    [1   :0]  s_1_axi_awburst;             
wire    [3   :0]  s_1_axi_awcache;             
wire    [7   :0]  s_1_axi_awid;                
wire    [7   :0]  s_1_axi_awlen;               
wire    [0   :0]  s_1_axi_awlock;              
wire    [2   :0]  s_1_axi_awprot;              
wire    [3   :0]  s_1_axi_awqos;               
wire              s_1_axi_awready;             
wire    [2   :0]  s_1_axi_awsize;              
wire              s_1_axi_awvalid;             
wire    [7   :0]  s_1_axi_bid;                 
wire              s_1_axi_bready;              
wire    [1   :0]  s_1_axi_bresp;               
wire              s_1_axi_bvalid;              
wire    [1023:0]  s_1_axi_rdata;               
wire    [7   :0]  s_1_axi_rid;                 
wire              s_1_axi_rlast;               
wire              s_1_axi_rready;              
wire    [1   :0]  s_1_axi_rresp;               
wire              s_1_axi_rvalid;              
wire    [1023:0]  s_1_axi_wdata;               
wire              s_1_axi_wlast;               
wire              s_1_axi_wready;              
wire    [127 :0]  s_1_axi_wstrb;               
wire              s_1_axi_wvalid;              
wire    [31  :0]  s_2_axi_araddr;              
wire    [1   :0]  s_2_axi_arburst;             
wire    [3   :0]  s_2_axi_arcache;             
wire    [7   :0]  s_2_axi_arid;                
wire    [7   :0]  s_2_axi_arlen;               
wire    [0   :0]  s_2_axi_arlock;              
wire    [2   :0]  s_2_axi_arprot;              
wire    [3   :0]  s_2_axi_arqos;               
wire              s_2_axi_arready;             
wire    [2   :0]  s_2_axi_arsize;              
wire              s_2_axi_arvalid;             
wire    [31  :0]  s_2_axi_awaddr;              
wire    [1   :0]  s_2_axi_awburst;             
wire    [3   :0]  s_2_axi_awcache;             
wire    [7   :0]  s_2_axi_awid;                
wire    [7   :0]  s_2_axi_awlen;               
wire    [0   :0]  s_2_axi_awlock;              
wire    [2   :0]  s_2_axi_awprot;              
wire    [3   :0]  s_2_axi_awqos;               
wire              s_2_axi_awready;             
wire    [2   :0]  s_2_axi_awsize;              
wire              s_2_axi_awvalid;             
wire    [7   :0]  s_2_axi_bid;                 
wire              s_2_axi_bready;              
wire    [1   :0]  s_2_axi_bresp;               
wire              s_2_axi_bvalid;              
wire    [1023:0]  s_2_axi_rdata;               
wire    [7   :0]  s_2_axi_rid;                 
wire              s_2_axi_rlast;               
wire              s_2_axi_rready;              
wire    [1   :0]  s_2_axi_rresp;               
wire              s_2_axi_rvalid;              
wire    [1023:0]  s_2_axi_wdata;               
wire              s_2_axi_wlast;               
wire              s_2_axi_wready;              
wire    [127 :0]  s_2_axi_wstrb;               
wire              s_2_axi_wvalid;              
wire    [31  :0]  s_3_axi_araddr;              
wire    [1   :0]  s_3_axi_arburst;             
wire    [3   :0]  s_3_axi_arcache;             
wire    [7   :0]  s_3_axi_arid;                
wire    [7   :0]  s_3_axi_arlen;               
wire    [0   :0]  s_3_axi_arlock;              
wire    [2   :0]  s_3_axi_arprot;              
wire    [3   :0]  s_3_axi_arqos;               
wire              s_3_axi_arready;             
wire    [2   :0]  s_3_axi_arsize;              
wire              s_3_axi_arvalid;             
wire    [31  :0]  s_3_axi_awaddr;              
wire    [1   :0]  s_3_axi_awburst;             
wire    [3   :0]  s_3_axi_awcache;             
wire    [7   :0]  s_3_axi_awid;                
wire    [7   :0]  s_3_axi_awlen;               
wire    [0   :0]  s_3_axi_awlock;              
wire    [2   :0]  s_3_axi_awprot;              
wire    [3   :0]  s_3_axi_awqos;               
wire              s_3_axi_awready;             
wire    [2   :0]  s_3_axi_awsize;              
wire              s_3_axi_awvalid;             
wire    [7   :0]  s_3_axi_bid;                 
wire              s_3_axi_bready;              
wire    [1   :0]  s_3_axi_bresp;               
wire              s_3_axi_bvalid;              
wire    [1023:0]  s_3_axi_rdata;               
wire    [7   :0]  s_3_axi_rid;                 
wire              s_3_axi_rlast;               
wire              s_3_axi_rready;              
wire    [1   :0]  s_3_axi_rresp;               
wire              s_3_axi_rvalid;              
wire    [1023:0]  s_3_axi_wdata;               
wire              s_3_axi_wlast;               
wire              s_3_axi_wready;              
wire    [127 :0]  s_3_axi_wstrb;               
wire              s_3_axi_wvalid;              


// Inst RV Cluster
// &Instance("rv_cluster_top"); @7
rv_cluster_top  x_rv_cluster_top (
  .rv_0_clk               (rv_0_clk              ),
  .rv_0_m_axi_araddr      (rv_0_m_axi_araddr     ),
  .rv_0_m_axi_arburst     (rv_0_m_axi_arburst    ),
  .rv_0_m_axi_arcache     (rv_0_m_axi_arcache    ),
  .rv_0_m_axi_arid        (rv_0_m_axi_arid       ),
  .rv_0_m_axi_arlen       (rv_0_m_axi_arlen      ),
  .rv_0_m_axi_arlock      (rv_0_m_axi_arlock     ),
  .rv_0_m_axi_arprot      (rv_0_m_axi_arprot     ),
  .rv_0_m_axi_arqos       (rv_0_m_axi_arqos      ),
  .rv_0_m_axi_arready     (rv_0_m_axi_arready    ),
  .rv_0_m_axi_arsize      (rv_0_m_axi_arsize     ),
  .rv_0_m_axi_arvalid     (rv_0_m_axi_arvalid    ),
  .rv_0_m_axi_awaddr      (rv_0_m_axi_awaddr     ),
  .rv_0_m_axi_awburst     (rv_0_m_axi_awburst    ),
  .rv_0_m_axi_awcache     (rv_0_m_axi_awcache    ),
  .rv_0_m_axi_awid        (rv_0_m_axi_awid       ),
  .rv_0_m_axi_awlen       (rv_0_m_axi_awlen      ),
  .rv_0_m_axi_awlock      (rv_0_m_axi_awlock     ),
  .rv_0_m_axi_awprot      (rv_0_m_axi_awprot     ),
  .rv_0_m_axi_awqos       (rv_0_m_axi_awqos      ),
  .rv_0_m_axi_awready     (rv_0_m_axi_awready    ),
  .rv_0_m_axi_awsize      (rv_0_m_axi_awsize     ),
  .rv_0_m_axi_awvalid     (rv_0_m_axi_awvalid    ),
  .rv_0_m_axi_bid         (rv_0_m_axi_bid        ),
  .rv_0_m_axi_bready      (rv_0_m_axi_bready     ),
  .rv_0_m_axi_bresp       (rv_0_m_axi_bresp      ),
  .rv_0_m_axi_bvalid      (rv_0_m_axi_bvalid     ),
  .rv_0_m_axi_rdata       (rv_0_m_axi_rdata      ),
  .rv_0_m_axi_rid         (rv_0_m_axi_rid        ),
  .rv_0_m_axi_rlast       (rv_0_m_axi_rlast      ),
  .rv_0_m_axi_rready      (rv_0_m_axi_rready     ),
  .rv_0_m_axi_rresp       (rv_0_m_axi_rresp      ),
  .rv_0_m_axi_rvalid      (rv_0_m_axi_rvalid     ),
  .rv_0_m_axi_wdata       (rv_0_m_axi_wdata      ),
  .rv_0_m_axi_wlast       (rv_0_m_axi_wlast      ),
  .rv_0_m_axi_wready      (rv_0_m_axi_wready     ),
  .rv_0_m_axi_wstrb       (rv_0_m_axi_wstrb      ),
  .rv_0_m_axi_wvalid      (rv_0_m_axi_wvalid     ),
  .rv_0_retire_pc         (rv_0_retire_pc        ),
  .rv_0_rst_addr          (rv_0_rst_addr         ),
  .rv_0_rstn              (rv_0_rstn             ),
  .rv_0_xocc_2_clk        (dsa_2_clk                   ),
  .rv_0_xocc_2_cmd_buffer (rv_0_xocc_2_cmd_buffer),
  .rv_0_xocc_2_cmd_empty  (rv_0_xocc_2_cmd_empty ),
  .rv_0_xocc_2_cmd_rd_en  (rv_0_xocc_2_cmd_rd_en ),
  .rv_0_xocc_2_rsp_buffer (rv_0_xocc_2_rsp_buffer),
  .rv_0_xocc_2_rsp_full   (rv_0_xocc_2_rsp_full  ),
  .rv_0_xocc_2_rsp_wr_en  (rv_0_xocc_2_rsp_wr_en ),
  .rv_0_xocc_2_rst        (dsa_2_rstn                  ),
  .rv_1_clk                (rv_1_clk               ),
  .rv_1_m_axi_araddr       (rv_1_m_axi_araddr      ),
  .rv_1_m_axi_arburst      (rv_1_m_axi_arburst     ),
  .rv_1_m_axi_arcache      (rv_1_m_axi_arcache     ),
  .rv_1_m_axi_arid         (rv_1_m_axi_arid        ),
  .rv_1_m_axi_arlen        (rv_1_m_axi_arlen       ),
  .rv_1_m_axi_arlock       (rv_1_m_axi_arlock      ),
  .rv_1_m_axi_arprot       (rv_1_m_axi_arprot      ),
  .rv_1_m_axi_arqos        (rv_1_m_axi_arqos       ),
  .rv_1_m_axi_arready      (rv_1_m_axi_arready     ),
  .rv_1_m_axi_arsize       (rv_1_m_axi_arsize      ),
  .rv_1_m_axi_arvalid      (rv_1_m_axi_arvalid     ),
  .rv_1_m_axi_awaddr       (rv_1_m_axi_awaddr      ),
  .rv_1_m_axi_awburst      (rv_1_m_axi_awburst     ),
  .rv_1_m_axi_awcache      (rv_1_m_axi_awcache     ),
  .rv_1_m_axi_awid         (rv_1_m_axi_awid        ),
  .rv_1_m_axi_awlen        (rv_1_m_axi_awlen       ),
  .rv_1_m_axi_awlock       (rv_1_m_axi_awlock      ),
  .rv_1_m_axi_awprot       (rv_1_m_axi_awprot      ),
  .rv_1_m_axi_awqos        (rv_1_m_axi_awqos       ),
  .rv_1_m_axi_awready      (rv_1_m_axi_awready     ),
  .rv_1_m_axi_awsize       (rv_1_m_axi_awsize      ),
  .rv_1_m_axi_awvalid      (rv_1_m_axi_awvalid     ),
  .rv_1_m_axi_bid          (rv_1_m_axi_bid         ),
  .rv_1_m_axi_bready       (rv_1_m_axi_bready      ),
  .rv_1_m_axi_bresp        (rv_1_m_axi_bresp       ),
  .rv_1_m_axi_bvalid       (rv_1_m_axi_bvalid      ),
  .rv_1_m_axi_rdata        (rv_1_m_axi_rdata       ),
  .rv_1_m_axi_rid          (rv_1_m_axi_rid         ),
  .rv_1_m_axi_rlast        (rv_1_m_axi_rlast       ),
  .rv_1_m_axi_rready       (rv_1_m_axi_rready      ),
  .rv_1_m_axi_rresp        (rv_1_m_axi_rresp       ),
  .rv_1_m_axi_rvalid       (rv_1_m_axi_rvalid      ),
  .rv_1_m_axi_wdata        (rv_1_m_axi_wdata       ),
  .rv_1_m_axi_wlast        (rv_1_m_axi_wlast       ),
  .rv_1_m_axi_wready       (rv_1_m_axi_wready      ),
  .rv_1_m_axi_wstrb        (rv_1_m_axi_wstrb       ),
  .rv_1_m_axi_wvalid       (rv_1_m_axi_wvalid      ),
  .rv_1_retire_pc          (rv_1_retire_pc         ),
  .rv_1_rst_addr           (rv_1_rst_addr          ),
  .rv_1_rstn               (rv_1_rstn              ),
  .rv_1_xocc_3_clk         (dsa_0_clk                   ),
  .rv_1_xocc_3_cmd_buffer  (rv_1_xocc_3_cmd_buffer ),
  .rv_1_xocc_3_cmd_empty   (rv_1_xocc_3_cmd_empty  ),
  .rv_1_xocc_3_cmd_rd_en   (rv_1_xocc_3_cmd_rd_en  ),
  .rv_1_xocc_3_rsp_buffer  (rv_1_xocc_3_rsp_buffer ),
  .rv_1_xocc_3_rsp_full    (rv_1_xocc_3_rsp_full   ),
  .rv_1_xocc_3_rsp_wr_en   (rv_1_xocc_3_rsp_wr_en  ),
  .rv_1_xocc_3_rst         (dsa_0_rstn                  ),
  .rv_2_clk                (rv_2_clk               ),
  .rv_2_m_axi_araddr       (rv_2_m_axi_araddr      ),
  .rv_2_m_axi_arburst      (rv_2_m_axi_arburst     ),
  .rv_2_m_axi_arcache      (rv_2_m_axi_arcache     ),
  .rv_2_m_axi_arid         (rv_2_m_axi_arid        ),
  .rv_2_m_axi_arlen        (rv_2_m_axi_arlen       ),
  .rv_2_m_axi_arlock       (rv_2_m_axi_arlock      ),
  .rv_2_m_axi_arprot       (rv_2_m_axi_arprot      ),
  .rv_2_m_axi_arqos        (rv_2_m_axi_arqos       ),
  .rv_2_m_axi_arready      (rv_2_m_axi_arready     ),
  .rv_2_m_axi_arsize       (rv_2_m_axi_arsize      ),
  .rv_2_m_axi_arvalid      (rv_2_m_axi_arvalid     ),
  .rv_2_m_axi_awaddr       (rv_2_m_axi_awaddr      ),
  .rv_2_m_axi_awburst      (rv_2_m_axi_awburst     ),
  .rv_2_m_axi_awcache      (rv_2_m_axi_awcache     ),
  .rv_2_m_axi_awid         (rv_2_m_axi_awid        ),
  .rv_2_m_axi_awlen        (rv_2_m_axi_awlen       ),
  .rv_2_m_axi_awlock       (rv_2_m_axi_awlock      ),
  .rv_2_m_axi_awprot       (rv_2_m_axi_awprot      ),
  .rv_2_m_axi_awqos        (rv_2_m_axi_awqos       ),
  .rv_2_m_axi_awready      (rv_2_m_axi_awready     ),
  .rv_2_m_axi_awsize       (rv_2_m_axi_awsize      ),
  .rv_2_m_axi_awvalid      (rv_2_m_axi_awvalid     ),
  .rv_2_m_axi_bid          (rv_2_m_axi_bid         ),
  .rv_2_m_axi_bready       (rv_2_m_axi_bready      ),
  .rv_2_m_axi_bresp        (rv_2_m_axi_bresp       ),
  .rv_2_m_axi_bvalid       (rv_2_m_axi_bvalid      ),
  .rv_2_m_axi_rdata        (rv_2_m_axi_rdata       ),
  .rv_2_m_axi_rid          (rv_2_m_axi_rid         ),
  .rv_2_m_axi_rlast        (rv_2_m_axi_rlast       ),
  .rv_2_m_axi_rready       (rv_2_m_axi_rready      ),
  .rv_2_m_axi_rresp        (rv_2_m_axi_rresp       ),
  .rv_2_m_axi_rvalid       (rv_2_m_axi_rvalid      ),
  .rv_2_m_axi_wdata        (rv_2_m_axi_wdata       ),
  .rv_2_m_axi_wlast        (rv_2_m_axi_wlast       ),
  .rv_2_m_axi_wready       (rv_2_m_axi_wready      ),
  .rv_2_m_axi_wstrb        (rv_2_m_axi_wstrb       ),
  .rv_2_m_axi_wvalid       (rv_2_m_axi_wvalid      ),
  .rv_2_retire_pc          (rv_2_retire_pc         ),
  .rv_2_rst_addr           (rv_2_rst_addr          ),
  .rv_2_rstn               (rv_2_rstn              ),
  .rv_2_xocc_4_clk         (dsa_1_clk                   ),
  .rv_2_xocc_4_cmd_buffer  (rv_2_xocc_4_cmd_buffer ),
  .rv_2_xocc_4_cmd_empty   (rv_2_xocc_4_cmd_empty  ),
  .rv_2_xocc_4_cmd_rd_en   (rv_2_xocc_4_cmd_rd_en  ),
  .rv_2_xocc_4_rsp_buffer  (rv_2_xocc_4_rsp_buffer ),
  .rv_2_xocc_4_rsp_full    (rv_2_xocc_4_rsp_full   ),
  .rv_2_xocc_4_rsp_wr_en   (rv_2_xocc_4_rsp_wr_en  ),
  .rv_2_xocc_4_rst         (dsa_1_rstn                  )
);

// &Connect( @8
//     .rv_0_xocc_2_clk (dsa_2_clk), @9
//     .rv_0_xocc_2_rst (dsa_2_rstn), @10
//     .rv_1_xocc_3_clk (dsa_0_clk), @11
//     .rv_1_xocc_3_rst (dsa_0_rstn), @12
//     .rv_2_xocc_4_clk (dsa_1_clk), @13
//     .rv_2_xocc_4_rst (dsa_1_rstn), @14
// ); @15

// Inst dsa_0 
// &ConnRule(s/dsa0_(\w+)_fifo/rv_1_xocc_3_$1/); @18
// &ConnRule(s/m00_axi/dsa_0_m_axi/); @19
// &Instance("dummy_dsa_wrapper", "x_dsa_0_top_wrapper"); @20
dummy_dsa_wrapper  x_dsa_0_top_wrapper (
  .clk                         (dsa_0_clk                  ),
  .dsa0_cmd_fifo_empty         (rv_1_xocc_3_cmd_empty ),
  .dsa0_cmd_fifo_rd_en         (rv_1_xocc_3_cmd_rd_en ),
  .dsa0_rsp_fifo_full          (rv_1_xocc_3_rsp_full  ),
  .dsa0_rsp_fifo_wr_en         (rv_1_xocc_3_rsp_wr_en ),
  .dsa0_xocc_cmd_in            (rv_1_xocc_3_cmd_buffer),
  .dsa0_xocc_cmd_out           (rv_1_xocc_3_rsp_buffer),
  .m00_axi_araddr              (dsa_0_m_axi_araddr         ),
  .m00_axi_arburst             (dsa_0_m_axi_arburst        ),
  .m00_axi_arcache             (dsa_0_m_axi_arcache        ),
  .m00_axi_arid                (dsa_0_m_axi_arid           ),
  .m00_axi_arlen               (dsa_0_m_axi_arlen          ),
  .m00_axi_arlock              (dsa_0_m_axi_arlock         ),
  .m00_axi_arprot              (dsa_0_m_axi_arprot         ),
  .m00_axi_arqos               (dsa_0_m_axi_arqos          ),
  .m00_axi_arready             (dsa_0_m_axi_arready        ),
  .m00_axi_arsize              (dsa_0_m_axi_arsize         ),
  .m00_axi_arvalid             (dsa_0_m_axi_arvalid        ),
  .m00_axi_awaddr              (dsa_0_m_axi_awaddr         ),
  .m00_axi_awburst             (dsa_0_m_axi_awburst        ),
  .m00_axi_awcache             (dsa_0_m_axi_awcache        ),
  .m00_axi_awid                (dsa_0_m_axi_awid           ),
  .m00_axi_awlen               (dsa_0_m_axi_awlen          ),
  .m00_axi_awlock              (dsa_0_m_axi_awlock         ),
  .m00_axi_awprot              (dsa_0_m_axi_awprot         ),
  .m00_axi_awqos               (dsa_0_m_axi_awqos          ),
  .m00_axi_awready             (dsa_0_m_axi_awready        ),
  .m00_axi_awsize              (dsa_0_m_axi_awsize         ),
  .m00_axi_awvalid             (dsa_0_m_axi_awvalid        ),
  .m00_axi_bid                 (dsa_0_m_axi_bid            ),
  .m00_axi_bready              (dsa_0_m_axi_bready         ),
  .m00_axi_bresp               (dsa_0_m_axi_bresp          ),
  .m00_axi_bvalid              (dsa_0_m_axi_bvalid         ),
  .m00_axi_rdata               (dsa_0_m_axi_rdata          ),
  .m00_axi_rid                 (dsa_0_m_axi_rid            ),
  .m00_axi_rlast               (dsa_0_m_axi_rlast          ),
  .m00_axi_rready              (dsa_0_m_axi_rready         ),
  .m00_axi_rresp               (dsa_0_m_axi_rresp          ),
  .m00_axi_rvalid              (dsa_0_m_axi_rvalid         ),
  .m00_axi_wdata               (dsa_0_m_axi_wdata          ),
  .m00_axi_wlast               (dsa_0_m_axi_wlast          ),
  .m00_axi_wready              (dsa_0_m_axi_wready         ),
  .m00_axi_wstrb               (dsa_0_m_axi_wstrb          ),
  .m00_axi_wvalid              (dsa_0_m_axi_wvalid         ),
  .rst                         (dsa_0_rstn                 )
);

// &Connect( @21
//     .dsa0_xocc_cmd_in (rv_1_xocc_3_cmd_buffer), @22
//     .dsa0_xocc_cmd_out(rv_1_xocc_3_rsp_buffer), @23
//     .clk(dsa_0_clk), @24
//     .rst(dsa_0_rstn), @25
// ); @26

// Inst dsa_1 
// &ConnRule(s/dsa0_(\w+)_fifo/rv_2_xocc_4_$1/); @29
// &ConnRule(s/m00_axi/dsa_1_m_axi/); @30
// &Instance("dummy_dsa_wrapper", "x_dsa_1_top_wrapper"); @31
dummy_dsa_wrapper  x_dsa_1_top_wrapper (
  .clk                         (dsa_1_clk                  ),
  .dsa0_cmd_fifo_empty         (rv_2_xocc_4_cmd_empty ),
  .dsa0_cmd_fifo_rd_en         (rv_2_xocc_4_cmd_rd_en ),
  .dsa0_rsp_fifo_full          (rv_2_xocc_4_rsp_full  ),
  .dsa0_rsp_fifo_wr_en         (rv_2_xocc_4_rsp_wr_en ),
  .dsa0_xocc_cmd_in            (rv_2_xocc_4_cmd_buffer),
  .dsa0_xocc_cmd_out           (rv_2_xocc_4_rsp_buffer),
  .m00_axi_araddr              (dsa_1_m_axi_araddr         ),
  .m00_axi_arburst             (dsa_1_m_axi_arburst        ),
  .m00_axi_arcache             (dsa_1_m_axi_arcache        ),
  .m00_axi_arid                (dsa_1_m_axi_arid           ),
  .m00_axi_arlen               (dsa_1_m_axi_arlen          ),
  .m00_axi_arlock              (dsa_1_m_axi_arlock         ),
  .m00_axi_arprot              (dsa_1_m_axi_arprot         ),
  .m00_axi_arqos               (dsa_1_m_axi_arqos          ),
  .m00_axi_arready             (dsa_1_m_axi_arready        ),
  .m00_axi_arsize              (dsa_1_m_axi_arsize         ),
  .m00_axi_arvalid             (dsa_1_m_axi_arvalid        ),
  .m00_axi_awaddr              (dsa_1_m_axi_awaddr         ),
  .m00_axi_awburst             (dsa_1_m_axi_awburst        ),
  .m00_axi_awcache             (dsa_1_m_axi_awcache        ),
  .m00_axi_awid                (dsa_1_m_axi_awid           ),
  .m00_axi_awlen               (dsa_1_m_axi_awlen          ),
  .m00_axi_awlock              (dsa_1_m_axi_awlock         ),
  .m00_axi_awprot              (dsa_1_m_axi_awprot         ),
  .m00_axi_awqos               (dsa_1_m_axi_awqos          ),
  .m00_axi_awready             (dsa_1_m_axi_awready        ),
  .m00_axi_awsize              (dsa_1_m_axi_awsize         ),
  .m00_axi_awvalid             (dsa_1_m_axi_awvalid        ),
  .m00_axi_bid                 (dsa_1_m_axi_bid            ),
  .m00_axi_bready              (dsa_1_m_axi_bready         ),
  .m00_axi_bresp               (dsa_1_m_axi_bresp          ),
  .m00_axi_bvalid              (dsa_1_m_axi_bvalid         ),
  .m00_axi_rdata               (dsa_1_m_axi_rdata          ),
  .m00_axi_rid                 (dsa_1_m_axi_rid            ),
  .m00_axi_rlast               (dsa_1_m_axi_rlast          ),
  .m00_axi_rready              (dsa_1_m_axi_rready         ),
  .m00_axi_rresp               (dsa_1_m_axi_rresp          ),
  .m00_axi_rvalid              (dsa_1_m_axi_rvalid         ),
  .m00_axi_wdata               (dsa_1_m_axi_wdata          ),
  .m00_axi_wlast               (dsa_1_m_axi_wlast          ),
  .m00_axi_wready              (dsa_1_m_axi_wready         ),
  .m00_axi_wstrb               (dsa_1_m_axi_wstrb          ),
  .m00_axi_wvalid              (dsa_1_m_axi_wvalid         ),
  .rst                         (dsa_1_rstn                 )
);

// &Connect( @32
//     .dsa0_xocc_cmd_in (rv_2_xocc_4_cmd_buffer), @33
//     .dsa0_xocc_cmd_out(rv_2_xocc_4_rsp_buffer), @34
//     .clk(dsa_1_clk), @35
//     .rst(dsa_1_rstn), @36
// ); @37

// Inst dsa_2 
// &ConnRule(s/dsa0_(\w+)_fifo/rv_0_xocc_2_$1/); @40
// &ConnRule(s/m00_axi/dsa_2_m_axi/); @41
// &Instance("dummy_dsa_wrapper", "x_dsa_2_top_wrapper"); @42
dummy_dsa_wrapper  x_dsa_2_top_wrapper (
  .clk                          (dsa_2_clk                   ),
  .dsa0_cmd_fifo_empty          (rv_0_xocc_2_cmd_empty ),
  .dsa0_cmd_fifo_rd_en          (rv_0_xocc_2_cmd_rd_en ),
  .dsa0_rsp_fifo_full           (rv_0_xocc_2_rsp_full  ),
  .dsa0_rsp_fifo_wr_en          (rv_0_xocc_2_rsp_wr_en ),
  .dsa0_xocc_cmd_in             (rv_0_xocc_2_cmd_buffer),
  .dsa0_xocc_cmd_out            (rv_0_xocc_2_rsp_buffer),
  .m00_axi_araddr               (dsa_2_m_axi_araddr          ),
  .m00_axi_arburst              (dsa_2_m_axi_arburst         ),
  .m00_axi_arcache              (dsa_2_m_axi_arcache         ),
  .m00_axi_arid                 (dsa_2_m_axi_arid            ),
  .m00_axi_arlen                (dsa_2_m_axi_arlen           ),
  .m00_axi_arlock               (dsa_2_m_axi_arlock          ),
  .m00_axi_arprot               (dsa_2_m_axi_arprot          ),
  .m00_axi_arqos                (dsa_2_m_axi_arqos           ),
  .m00_axi_arready              (dsa_2_m_axi_arready         ),
  .m00_axi_arsize               (dsa_2_m_axi_arsize          ),
  .m00_axi_arvalid              (dsa_2_m_axi_arvalid         ),
  .m00_axi_awaddr               (dsa_2_m_axi_awaddr          ),
  .m00_axi_awburst              (dsa_2_m_axi_awburst         ),
  .m00_axi_awcache              (dsa_2_m_axi_awcache         ),
  .m00_axi_awid                 (dsa_2_m_axi_awid            ),
  .m00_axi_awlen                (dsa_2_m_axi_awlen           ),
  .m00_axi_awlock               (dsa_2_m_axi_awlock          ),
  .m00_axi_awprot               (dsa_2_m_axi_awprot          ),
  .m00_axi_awqos                (dsa_2_m_axi_awqos           ),
  .m00_axi_awready              (dsa_2_m_axi_awready         ),
  .m00_axi_awsize               (dsa_2_m_axi_awsize          ),
  .m00_axi_awvalid              (dsa_2_m_axi_awvalid         ),
  .m00_axi_bid                  (dsa_2_m_axi_bid             ),
  .m00_axi_bready               (dsa_2_m_axi_bready          ),
  .m00_axi_bresp                (dsa_2_m_axi_bresp           ),
  .m00_axi_bvalid               (dsa_2_m_axi_bvalid          ),
  .m00_axi_rdata                (dsa_2_m_axi_rdata           ),
  .m00_axi_rid                  (dsa_2_m_axi_rid             ),
  .m00_axi_rlast                (dsa_2_m_axi_rlast           ),
  .m00_axi_rready               (dsa_2_m_axi_rready          ),
  .m00_axi_rresp                (dsa_2_m_axi_rresp           ),
  .m00_axi_rvalid               (dsa_2_m_axi_rvalid          ),
  .m00_axi_wdata                (dsa_2_m_axi_wdata           ),
  .m00_axi_wlast                (dsa_2_m_axi_wlast           ),
  .m00_axi_wready               (dsa_2_m_axi_wready          ),
  .m00_axi_wstrb                (dsa_2_m_axi_wstrb           ),
  .m00_axi_wvalid               (dsa_2_m_axi_wvalid          ),
  .rst                          (dsa_2_rstn                  )
);

// &Connect( @43
//     .dsa0_xocc_cmd_in (rv_0_xocc_2_cmd_buffer), @44
//     .dsa0_xocc_cmd_out(rv_0_xocc_2_rsp_buffer), @45
//     .clk(dsa_2_clk), @46
//     .rst(dsa_2_rstn), @47
// ); @48

// Mem SS
// &Instance("mem_sub_sys_top"); @51
mem_sub_sys_top  x_mem_sub_sys_top (
  .mem_sub_sys_clk  (mem_sub_sys_clk ),
  .mem_sub_sys_rstn (mem_sub_sys_rstn),
  .s_0_axi_araddr   (s_0_axi_araddr  ),
  .s_0_axi_arburst  (s_0_axi_arburst ),
  .s_0_axi_arcache  (s_0_axi_arcache ),
  .s_0_axi_arid     (s_0_axi_arid    ),
  .s_0_axi_arlen    (s_0_axi_arlen   ),
  .s_0_axi_arlock   (s_0_axi_arlock  ),
  .s_0_axi_arprot   (s_0_axi_arprot  ),
  .s_0_axi_arqos    (s_0_axi_arqos   ),
  .s_0_axi_arready  (s_0_axi_arready ),
  .s_0_axi_arsize   (s_0_axi_arsize  ),
  .s_0_axi_arvalid  (s_0_axi_arvalid ),
  .s_0_axi_awaddr   (s_0_axi_awaddr  ),
  .s_0_axi_awburst  (s_0_axi_awburst ),
  .s_0_axi_awcache  (s_0_axi_awcache ),
  .s_0_axi_awid     (s_0_axi_awid    ),
  .s_0_axi_awlen    (s_0_axi_awlen   ),
  .s_0_axi_awlock   (s_0_axi_awlock  ),
  .s_0_axi_awprot   (s_0_axi_awprot  ),
  .s_0_axi_awqos    (s_0_axi_awqos   ),
  .s_0_axi_awready  (s_0_axi_awready ),
  .s_0_axi_awsize   (s_0_axi_awsize  ),
  .s_0_axi_awvalid  (s_0_axi_awvalid ),
  .s_0_axi_bid      (s_0_axi_bid     ),
  .s_0_axi_bready   (s_0_axi_bready  ),
  .s_0_axi_bresp    (s_0_axi_bresp   ),
  .s_0_axi_bvalid   (s_0_axi_bvalid  ),
  .s_0_axi_rdata    (s_0_axi_rdata   ),
  .s_0_axi_rid      (s_0_axi_rid     ),
  .s_0_axi_rlast    (s_0_axi_rlast   ),
  .s_0_axi_rready   (s_0_axi_rready  ),
  .s_0_axi_rresp    (s_0_axi_rresp   ),
  .s_0_axi_rvalid   (s_0_axi_rvalid  ),
  .s_0_axi_wdata    (s_0_axi_wdata   ),
  .s_0_axi_wlast    (s_0_axi_wlast   ),
  .s_0_axi_wready   (s_0_axi_wready  ),
  .s_0_axi_wstrb    (s_0_axi_wstrb   ),
  .s_0_axi_wvalid   (s_0_axi_wvalid  ),
  .s_1_axi_araddr   (s_1_axi_araddr  ),
  .s_1_axi_arburst  (s_1_axi_arburst ),
  .s_1_axi_arcache  (s_1_axi_arcache ),
  .s_1_axi_arid     (s_1_axi_arid    ),
  .s_1_axi_arlen    (s_1_axi_arlen   ),
  .s_1_axi_arlock   (s_1_axi_arlock  ),
  .s_1_axi_arprot   (s_1_axi_arprot  ),
  .s_1_axi_arqos    (s_1_axi_arqos   ),
  .s_1_axi_arready  (s_1_axi_arready ),
  .s_1_axi_arsize   (s_1_axi_arsize  ),
  .s_1_axi_arvalid  (s_1_axi_arvalid ),
  .s_1_axi_awaddr   (s_1_axi_awaddr  ),
  .s_1_axi_awburst  (s_1_axi_awburst ),
  .s_1_axi_awcache  (s_1_axi_awcache ),
  .s_1_axi_awid     (s_1_axi_awid    ),
  .s_1_axi_awlen    (s_1_axi_awlen   ),
  .s_1_axi_awlock   (s_1_axi_awlock  ),
  .s_1_axi_awprot   (s_1_axi_awprot  ),
  .s_1_axi_awqos    (s_1_axi_awqos   ),
  .s_1_axi_awready  (s_1_axi_awready ),
  .s_1_axi_awsize   (s_1_axi_awsize  ),
  .s_1_axi_awvalid  (s_1_axi_awvalid ),
  .s_1_axi_bid      (s_1_axi_bid     ),
  .s_1_axi_bready   (s_1_axi_bready  ),
  .s_1_axi_bresp    (s_1_axi_bresp   ),
  .s_1_axi_bvalid   (s_1_axi_bvalid  ),
  .s_1_axi_rdata    (s_1_axi_rdata   ),
  .s_1_axi_rid      (s_1_axi_rid     ),
  .s_1_axi_rlast    (s_1_axi_rlast   ),
  .s_1_axi_rready   (s_1_axi_rready  ),
  .s_1_axi_rresp    (s_1_axi_rresp   ),
  .s_1_axi_rvalid   (s_1_axi_rvalid  ),
  .s_1_axi_wdata    (s_1_axi_wdata   ),
  .s_1_axi_wlast    (s_1_axi_wlast   ),
  .s_1_axi_wready   (s_1_axi_wready  ),
  .s_1_axi_wstrb    (s_1_axi_wstrb   ),
  .s_1_axi_wvalid   (s_1_axi_wvalid  ),
  .s_2_axi_araddr   (s_2_axi_araddr  ),
  .s_2_axi_arburst  (s_2_axi_arburst ),
  .s_2_axi_arcache  (s_2_axi_arcache ),
  .s_2_axi_arid     (s_2_axi_arid    ),
  .s_2_axi_arlen    (s_2_axi_arlen   ),
  .s_2_axi_arlock   (s_2_axi_arlock  ),
  .s_2_axi_arprot   (s_2_axi_arprot  ),
  .s_2_axi_arqos    (s_2_axi_arqos   ),
  .s_2_axi_arready  (s_2_axi_arready ),
  .s_2_axi_arsize   (s_2_axi_arsize  ),
  .s_2_axi_arvalid  (s_2_axi_arvalid ),
  .s_2_axi_awaddr   (s_2_axi_awaddr  ),
  .s_2_axi_awburst  (s_2_axi_awburst ),
  .s_2_axi_awcache  (s_2_axi_awcache ),
  .s_2_axi_awid     (s_2_axi_awid    ),
  .s_2_axi_awlen    (s_2_axi_awlen   ),
  .s_2_axi_awlock   (s_2_axi_awlock  ),
  .s_2_axi_awprot   (s_2_axi_awprot  ),
  .s_2_axi_awqos    (s_2_axi_awqos   ),
  .s_2_axi_awready  (s_2_axi_awready ),
  .s_2_axi_awsize   (s_2_axi_awsize  ),
  .s_2_axi_awvalid  (s_2_axi_awvalid ),
  .s_2_axi_bid      (s_2_axi_bid     ),
  .s_2_axi_bready   (s_2_axi_bready  ),
  .s_2_axi_bresp    (s_2_axi_bresp   ),
  .s_2_axi_bvalid   (s_2_axi_bvalid  ),
  .s_2_axi_rdata    (s_2_axi_rdata   ),
  .s_2_axi_rid      (s_2_axi_rid     ),
  .s_2_axi_rlast    (s_2_axi_rlast   ),
  .s_2_axi_rready   (s_2_axi_rready  ),
  .s_2_axi_rresp    (s_2_axi_rresp   ),
  .s_2_axi_rvalid   (s_2_axi_rvalid  ),
  .s_2_axi_wdata    (s_2_axi_wdata   ),
  .s_2_axi_wlast    (s_2_axi_wlast   ),
  .s_2_axi_wready   (s_2_axi_wready  ),
  .s_2_axi_wstrb    (s_2_axi_wstrb   ),
  .s_2_axi_wvalid   (s_2_axi_wvalid  ),
  .s_3_axi_araddr   (s_3_axi_araddr  ),
  .s_3_axi_arburst  (s_3_axi_arburst ),
  .s_3_axi_arcache  (s_3_axi_arcache ),
  .s_3_axi_arid     (s_3_axi_arid    ),
  .s_3_axi_arlen    (s_3_axi_arlen   ),
  .s_3_axi_arlock   (s_3_axi_arlock  ),
  .s_3_axi_arprot   (s_3_axi_arprot  ),
  .s_3_axi_arqos    (s_3_axi_arqos   ),
  .s_3_axi_arready  (s_3_axi_arready ),
  .s_3_axi_arsize   (s_3_axi_arsize  ),
  .s_3_axi_arvalid  (s_3_axi_arvalid ),
  .s_3_axi_awaddr   (s_3_axi_awaddr  ),
  .s_3_axi_awburst  (s_3_axi_awburst ),
  .s_3_axi_awcache  (s_3_axi_awcache ),
  .s_3_axi_awid     (s_3_axi_awid    ),
  .s_3_axi_awlen    (s_3_axi_awlen   ),
  .s_3_axi_awlock   (s_3_axi_awlock  ),
  .s_3_axi_awprot   (s_3_axi_awprot  ),
  .s_3_axi_awqos    (s_3_axi_awqos   ),
  .s_3_axi_awready  (s_3_axi_awready ),
  .s_3_axi_awsize   (s_3_axi_awsize  ),
  .s_3_axi_awvalid  (s_3_axi_awvalid ),
  .s_3_axi_bid      (s_3_axi_bid     ),
  .s_3_axi_bready   (s_3_axi_bready  ),
  .s_3_axi_bresp    (s_3_axi_bresp   ),
  .s_3_axi_bvalid   (s_3_axi_bvalid  ),
  .s_3_axi_rdata    (s_3_axi_rdata   ),
  .s_3_axi_rid      (s_3_axi_rid     ),
  .s_3_axi_rlast    (s_3_axi_rlast   ),
  .s_3_axi_rready   (s_3_axi_rready  ),
  .s_3_axi_rresp    (s_3_axi_rresp   ),
  .s_3_axi_rvalid   (s_3_axi_rvalid  ),
  .s_3_axi_wdata    (s_3_axi_wdata   ),
  .s_3_axi_wlast    (s_3_axi_wlast   ),
  .s_3_axi_wready   (s_3_axi_wready  ),
  .s_3_axi_wstrb    (s_3_axi_wstrb   ),
  .s_3_axi_wvalid   (s_3_axi_wvalid  )
);


// XBar
// &ConnRule(s/S00_AXI/rv_0_m_axi/); @54
// &ConnRule(s/S01_AXI/rv_1_m_axi/); @55
// &ConnRule(s/S02_AXI/rv_2_m_axi/); @56
// &ConnRule(s/S03_AXI/dsa_0_m_axi/); @57
// &ConnRule(s/S04_AXI/dsa_1_m_axi/); @58
// &ConnRule(s/S05_AXI/dsa_2_m_axi/); @59
// &ConnRule(s/M00_AXI/s_0_axi/); @60
// &ConnRule(s/M01_AXI/s_1_axi/); @61
// &ConnRule(s/M02_AXI/s_2_axi/); @62
// &ConnRule(s/M03_AXI/s_3_axi/); @63
// &Instance("xbar_top_wrapper"); @64
xbar_top_wrapper  x_xbar_top_wrapper (
  .M00_AXI_aclk             (mem_sub_sys_clk         ),
  .M00_AXI_araddr           (s_0_axi_araddr          ),
  .M00_AXI_arburst          (s_0_axi_arburst         ),
  .M00_AXI_arcache          (s_0_axi_arcache         ),
  .M00_AXI_aresetn          (mem_sub_sys_rstn        ),
  .M00_AXI_arid             (s_0_axi_arid            ),
  .M00_AXI_arlen            (s_0_axi_arlen           ),
  .M00_AXI_arlock           (s_0_axi_arlock          ),
  .M00_AXI_arprot           (s_0_axi_arprot          ),
  .M00_AXI_arqos            (s_0_axi_arqos           ),
  .M00_AXI_arready          (s_0_axi_arready         ),
  .M00_AXI_arsize           (s_0_axi_arsize          ),
  .M00_AXI_arvalid          (s_0_axi_arvalid         ),
  .M00_AXI_awaddr           (s_0_axi_awaddr          ),
  .M00_AXI_awburst          (s_0_axi_awburst         ),
  .M00_AXI_awcache          (s_0_axi_awcache         ),
  .M00_AXI_awid             (s_0_axi_awid            ),
  .M00_AXI_awlen            (s_0_axi_awlen           ),
  .M00_AXI_awlock           (s_0_axi_awlock          ),
  .M00_AXI_awprot           (s_0_axi_awprot          ),
  .M00_AXI_awqos            (s_0_axi_awqos           ),
  .M00_AXI_awready          (s_0_axi_awready         ),
  .M00_AXI_awsize           (s_0_axi_awsize          ),
  .M00_AXI_awvalid          (s_0_axi_awvalid         ),
  .M00_AXI_bid              (s_0_axi_bid             ),
  .M00_AXI_bready           (s_0_axi_bready          ),
  .M00_AXI_bresp            (s_0_axi_bresp           ),
  .M00_AXI_bvalid           (s_0_axi_bvalid          ),
  .M00_AXI_rdata            (s_0_axi_rdata           ),
  .M00_AXI_rid              (s_0_axi_rid             ),
  .M00_AXI_rlast            (s_0_axi_rlast           ),
  .M00_AXI_rready           (s_0_axi_rready          ),
  .M00_AXI_rresp            (s_0_axi_rresp           ),
  .M00_AXI_rvalid           (s_0_axi_rvalid          ),
  .M00_AXI_wdata            (s_0_axi_wdata           ),
  .M00_AXI_wlast            (s_0_axi_wlast           ),
  .M00_AXI_wready           (s_0_axi_wready          ),
  .M00_AXI_wstrb            (s_0_axi_wstrb           ),
  .M00_AXI_wvalid           (s_0_axi_wvalid          ),
  .M01_AXI_aclk             (mem_sub_sys_clk         ),
  .M01_AXI_araddr           (s_1_axi_araddr          ),
  .M01_AXI_arburst          (s_1_axi_arburst         ),
  .M01_AXI_arcache          (s_1_axi_arcache         ),
  .M01_AXI_aresetn          (mem_sub_sys_rstn        ),
  .M01_AXI_arid             (s_1_axi_arid            ),
  .M01_AXI_arlen            (s_1_axi_arlen           ),
  .M01_AXI_arlock           (s_1_axi_arlock          ),
  .M01_AXI_arprot           (s_1_axi_arprot          ),
  .M01_AXI_arqos            (s_1_axi_arqos           ),
  .M01_AXI_arready          (s_1_axi_arready         ),
  .M01_AXI_arsize           (s_1_axi_arsize          ),
  .M01_AXI_arvalid          (s_1_axi_arvalid         ),
  .M01_AXI_awaddr           (s_1_axi_awaddr          ),
  .M01_AXI_awburst          (s_1_axi_awburst         ),
  .M01_AXI_awcache          (s_1_axi_awcache         ),
  .M01_AXI_awid             (s_1_axi_awid            ),
  .M01_AXI_awlen            (s_1_axi_awlen           ),
  .M01_AXI_awlock           (s_1_axi_awlock          ),
  .M01_AXI_awprot           (s_1_axi_awprot          ),
  .M01_AXI_awqos            (s_1_axi_awqos           ),
  .M01_AXI_awready          (s_1_axi_awready         ),
  .M01_AXI_awsize           (s_1_axi_awsize          ),
  .M01_AXI_awvalid          (s_1_axi_awvalid         ),
  .M01_AXI_bid              (s_1_axi_bid             ),
  .M01_AXI_bready           (s_1_axi_bready          ),
  .M01_AXI_bresp            (s_1_axi_bresp           ),
  .M01_AXI_bvalid           (s_1_axi_bvalid          ),
  .M01_AXI_rdata            (s_1_axi_rdata           ),
  .M01_AXI_rid              (s_1_axi_rid             ),
  .M01_AXI_rlast            (s_1_axi_rlast           ),
  .M01_AXI_rready           (s_1_axi_rready          ),
  .M01_AXI_rresp            (s_1_axi_rresp           ),
  .M01_AXI_rvalid           (s_1_axi_rvalid          ),
  .M01_AXI_wdata            (s_1_axi_wdata           ),
  .M01_AXI_wlast            (s_1_axi_wlast           ),
  .M01_AXI_wready           (s_1_axi_wready          ),
  .M01_AXI_wstrb            (s_1_axi_wstrb           ),
  .M01_AXI_wvalid           (s_1_axi_wvalid          ),
  .M02_AXI_aclk             (mem_sub_sys_clk         ),
  .M02_AXI_araddr           (s_2_axi_araddr          ),
  .M02_AXI_arburst          (s_2_axi_arburst         ),
  .M02_AXI_arcache          (s_2_axi_arcache         ),
  .M02_AXI_aresetn          (mem_sub_sys_rstn        ),
  .M02_AXI_arid             (s_2_axi_arid            ),
  .M02_AXI_arlen            (s_2_axi_arlen           ),
  .M02_AXI_arlock           (s_2_axi_arlock          ),
  .M02_AXI_arprot           (s_2_axi_arprot          ),
  .M02_AXI_arqos            (s_2_axi_arqos           ),
  .M02_AXI_arready          (s_2_axi_arready         ),
  .M02_AXI_arsize           (s_2_axi_arsize          ),
  .M02_AXI_arvalid          (s_2_axi_arvalid         ),
  .M02_AXI_awaddr           (s_2_axi_awaddr          ),
  .M02_AXI_awburst          (s_2_axi_awburst         ),
  .M02_AXI_awcache          (s_2_axi_awcache         ),
  .M02_AXI_awid             (s_2_axi_awid            ),
  .M02_AXI_awlen            (s_2_axi_awlen           ),
  .M02_AXI_awlock           (s_2_axi_awlock          ),
  .M02_AXI_awprot           (s_2_axi_awprot          ),
  .M02_AXI_awqos            (s_2_axi_awqos           ),
  .M02_AXI_awready          (s_2_axi_awready         ),
  .M02_AXI_awsize           (s_2_axi_awsize          ),
  .M02_AXI_awvalid          (s_2_axi_awvalid         ),
  .M02_AXI_bid              (s_2_axi_bid             ),
  .M02_AXI_bready           (s_2_axi_bready          ),
  .M02_AXI_bresp            (s_2_axi_bresp           ),
  .M02_AXI_bvalid           (s_2_axi_bvalid          ),
  .M02_AXI_rdata            (s_2_axi_rdata           ),
  .M02_AXI_rid              (s_2_axi_rid             ),
  .M02_AXI_rlast            (s_2_axi_rlast           ),
  .M02_AXI_rready           (s_2_axi_rready          ),
  .M02_AXI_rresp            (s_2_axi_rresp           ),
  .M02_AXI_rvalid           (s_2_axi_rvalid          ),
  .M02_AXI_wdata            (s_2_axi_wdata           ),
  .M02_AXI_wlast            (s_2_axi_wlast           ),
  .M02_AXI_wready           (s_2_axi_wready          ),
  .M02_AXI_wstrb            (s_2_axi_wstrb           ),
  .M02_AXI_wvalid           (s_2_axi_wvalid          ),
  .M03_AXI_aclk             (mem_sub_sys_clk         ),
  .M03_AXI_araddr           (s_3_axi_araddr          ),
  .M03_AXI_arburst          (s_3_axi_arburst         ),
  .M03_AXI_arcache          (s_3_axi_arcache         ),
  .M03_AXI_aresetn          (mem_sub_sys_rstn        ),
  .M03_AXI_arid             (s_3_axi_arid            ),
  .M03_AXI_arlen            (s_3_axi_arlen           ),
  .M03_AXI_arlock           (s_3_axi_arlock          ),
  .M03_AXI_arprot           (s_3_axi_arprot          ),
  .M03_AXI_arqos            (s_3_axi_arqos           ),
  .M03_AXI_arready          (s_3_axi_arready         ),
  .M03_AXI_arsize           (s_3_axi_arsize          ),
  .M03_AXI_arvalid          (s_3_axi_arvalid         ),
  .M03_AXI_awaddr           (s_3_axi_awaddr          ),
  .M03_AXI_awburst          (s_3_axi_awburst         ),
  .M03_AXI_awcache          (s_3_axi_awcache         ),
  .M03_AXI_awid             (s_3_axi_awid            ),
  .M03_AXI_awlen            (s_3_axi_awlen           ),
  .M03_AXI_awlock           (s_3_axi_awlock          ),
  .M03_AXI_awprot           (s_3_axi_awprot          ),
  .M03_AXI_awqos            (s_3_axi_awqos           ),
  .M03_AXI_awready          (s_3_axi_awready         ),
  .M03_AXI_awsize           (s_3_axi_awsize          ),
  .M03_AXI_awvalid          (s_3_axi_awvalid         ),
  .M03_AXI_bid              (s_3_axi_bid             ),
  .M03_AXI_bready           (s_3_axi_bready          ),
  .M03_AXI_bresp            (s_3_axi_bresp           ),
  .M03_AXI_bvalid           (s_3_axi_bvalid          ),
  .M03_AXI_rdata            (s_3_axi_rdata           ),
  .M03_AXI_rid              (s_3_axi_rid             ),
  .M03_AXI_rlast            (s_3_axi_rlast           ),
  .M03_AXI_rready           (s_3_axi_rready          ),
  .M03_AXI_rresp            (s_3_axi_rresp           ),
  .M03_AXI_rvalid           (s_3_axi_rvalid          ),
  .M03_AXI_wdata            (s_3_axi_wdata           ),
  .M03_AXI_wlast            (s_3_axi_wlast           ),
  .M03_AXI_wready           (s_3_axi_wready          ),
  .M03_AXI_wstrb            (s_3_axi_wstrb           ),
  .M03_AXI_wvalid           (s_3_axi_wvalid          ),
  .S00_AXI_aclk             (rv_0_clk          ),
  .S00_AXI_araddr           (rv_0_m_axi_araddr ),
  .S00_AXI_arburst          (rv_0_m_axi_arburst),
  .S00_AXI_arcache          (rv_0_m_axi_arcache),
  .S00_AXI_aresetn          (rv_0_rstn         ),
  .S00_AXI_arid             (rv_0_m_axi_arid   ),
  .S00_AXI_arlen            (rv_0_m_axi_arlen  ),
  .S00_AXI_arlock           (rv_0_m_axi_arlock ),
  .S00_AXI_arprot           (rv_0_m_axi_arprot ),
  .S00_AXI_arqos            (rv_0_m_axi_arqos  ),
  .S00_AXI_arready          (rv_0_m_axi_arready),
  .S00_AXI_arsize           (rv_0_m_axi_arsize ),
  .S00_AXI_arvalid          (rv_0_m_axi_arvalid),
  .S00_AXI_awaddr           (rv_0_m_axi_awaddr ),
  .S00_AXI_awburst          (rv_0_m_axi_awburst),
  .S00_AXI_awcache          (rv_0_m_axi_awcache),
  .S00_AXI_awid             (rv_0_m_axi_awid   ),
  .S00_AXI_awlen            (rv_0_m_axi_awlen  ),
  .S00_AXI_awlock           (rv_0_m_axi_awlock ),
  .S00_AXI_awprot           (rv_0_m_axi_awprot ),
  .S00_AXI_awqos            (rv_0_m_axi_awqos  ),
  .S00_AXI_awready          (rv_0_m_axi_awready),
  .S00_AXI_awsize           (rv_0_m_axi_awsize ),
  .S00_AXI_awvalid          (rv_0_m_axi_awvalid),
  .S00_AXI_bid              (rv_0_m_axi_bid    ),
  .S00_AXI_bready           (rv_0_m_axi_bready ),
  .S00_AXI_bresp            (rv_0_m_axi_bresp  ),
  .S00_AXI_bvalid           (rv_0_m_axi_bvalid ),
  .S00_AXI_rdata            (rv_0_m_axi_rdata  ),
  .S00_AXI_rid              (rv_0_m_axi_rid    ),
  .S00_AXI_rlast            (rv_0_m_axi_rlast  ),
  .S00_AXI_rready           (rv_0_m_axi_rready ),
  .S00_AXI_rresp            (rv_0_m_axi_rresp  ),
  .S00_AXI_rvalid           (rv_0_m_axi_rvalid ),
  .S00_AXI_wdata            (rv_0_m_axi_wdata  ),
  .S00_AXI_wlast            (rv_0_m_axi_wlast  ),
  .S00_AXI_wready           (rv_0_m_axi_wready ),
  .S00_AXI_wstrb            (rv_0_m_axi_wstrb  ),
  .S00_AXI_wvalid           (rv_0_m_axi_wvalid ),
  .S01_AXI_aclk             (rv_1_clk           ),
  .S01_AXI_araddr           (rv_1_m_axi_araddr  ),
  .S01_AXI_arburst          (rv_1_m_axi_arburst ),
  .S01_AXI_arcache          (rv_1_m_axi_arcache ),
  .S01_AXI_aresetn          (rv_1_rstn          ),
  .S01_AXI_arid             (rv_1_m_axi_arid    ),
  .S01_AXI_arlen            (rv_1_m_axi_arlen   ),
  .S01_AXI_arlock           (rv_1_m_axi_arlock  ),
  .S01_AXI_arprot           (rv_1_m_axi_arprot  ),
  .S01_AXI_arqos            (rv_1_m_axi_arqos   ),
  .S01_AXI_arready          (rv_1_m_axi_arready ),
  .S01_AXI_arsize           (rv_1_m_axi_arsize  ),
  .S01_AXI_arvalid          (rv_1_m_axi_arvalid ),
  .S01_AXI_awaddr           (rv_1_m_axi_awaddr  ),
  .S01_AXI_awburst          (rv_1_m_axi_awburst ),
  .S01_AXI_awcache          (rv_1_m_axi_awcache ),
  .S01_AXI_awid             (rv_1_m_axi_awid    ),
  .S01_AXI_awlen            (rv_1_m_axi_awlen   ),
  .S01_AXI_awlock           (rv_1_m_axi_awlock  ),
  .S01_AXI_awprot           (rv_1_m_axi_awprot  ),
  .S01_AXI_awqos            (rv_1_m_axi_awqos   ),
  .S01_AXI_awready          (rv_1_m_axi_awready ),
  .S01_AXI_awsize           (rv_1_m_axi_awsize  ),
  .S01_AXI_awvalid          (rv_1_m_axi_awvalid ),
  .S01_AXI_bid              (rv_1_m_axi_bid     ),
  .S01_AXI_bready           (rv_1_m_axi_bready  ),
  .S01_AXI_bresp            (rv_1_m_axi_bresp   ),
  .S01_AXI_bvalid           (rv_1_m_axi_bvalid  ),
  .S01_AXI_rdata            (rv_1_m_axi_rdata   ),
  .S01_AXI_rid              (rv_1_m_axi_rid     ),
  .S01_AXI_rlast            (rv_1_m_axi_rlast   ),
  .S01_AXI_rready           (rv_1_m_axi_rready  ),
  .S01_AXI_rresp            (rv_1_m_axi_rresp   ),
  .S01_AXI_rvalid           (rv_1_m_axi_rvalid  ),
  .S01_AXI_wdata            (rv_1_m_axi_wdata   ),
  .S01_AXI_wlast            (rv_1_m_axi_wlast   ),
  .S01_AXI_wready           (rv_1_m_axi_wready  ),
  .S01_AXI_wstrb            (rv_1_m_axi_wstrb   ),
  .S01_AXI_wvalid           (rv_1_m_axi_wvalid  ),
  .S02_AXI_aclk             (rv_2_clk           ),
  .S02_AXI_araddr           (rv_2_m_axi_araddr  ),
  .S02_AXI_arburst          (rv_2_m_axi_arburst ),
  .S02_AXI_arcache          (rv_2_m_axi_arcache ),
  .S02_AXI_aresetn          (rv_2_rstn          ),
  .S02_AXI_arid             (rv_2_m_axi_arid    ),
  .S02_AXI_arlen            (rv_2_m_axi_arlen   ),
  .S02_AXI_arlock           (rv_2_m_axi_arlock  ),
  .S02_AXI_arprot           (rv_2_m_axi_arprot  ),
  .S02_AXI_arqos            (rv_2_m_axi_arqos   ),
  .S02_AXI_arready          (rv_2_m_axi_arready ),
  .S02_AXI_arsize           (rv_2_m_axi_arsize  ),
  .S02_AXI_arvalid          (rv_2_m_axi_arvalid ),
  .S02_AXI_awaddr           (rv_2_m_axi_awaddr  ),
  .S02_AXI_awburst          (rv_2_m_axi_awburst ),
  .S02_AXI_awcache          (rv_2_m_axi_awcache ),
  .S02_AXI_awid             (rv_2_m_axi_awid    ),
  .S02_AXI_awlen            (rv_2_m_axi_awlen   ),
  .S02_AXI_awlock           (rv_2_m_axi_awlock  ),
  .S02_AXI_awprot           (rv_2_m_axi_awprot  ),
  .S02_AXI_awqos            (rv_2_m_axi_awqos   ),
  .S02_AXI_awready          (rv_2_m_axi_awready ),
  .S02_AXI_awsize           (rv_2_m_axi_awsize  ),
  .S02_AXI_awvalid          (rv_2_m_axi_awvalid ),
  .S02_AXI_bid              (rv_2_m_axi_bid     ),
  .S02_AXI_bready           (rv_2_m_axi_bready  ),
  .S02_AXI_bresp            (rv_2_m_axi_bresp   ),
  .S02_AXI_bvalid           (rv_2_m_axi_bvalid  ),
  .S02_AXI_rdata            (rv_2_m_axi_rdata   ),
  .S02_AXI_rid              (rv_2_m_axi_rid     ),
  .S02_AXI_rlast            (rv_2_m_axi_rlast   ),
  .S02_AXI_rready           (rv_2_m_axi_rready  ),
  .S02_AXI_rresp            (rv_2_m_axi_rresp   ),
  .S02_AXI_rvalid           (rv_2_m_axi_rvalid  ),
  .S02_AXI_wdata            (rv_2_m_axi_wdata   ),
  .S02_AXI_wlast            (rv_2_m_axi_wlast   ),
  .S02_AXI_wready           (rv_2_m_axi_wready  ),
  .S02_AXI_wstrb            (rv_2_m_axi_wstrb   ),
  .S02_AXI_wvalid           (rv_2_m_axi_wvalid  ),
  .S03_AXI_aclk             (dsa_0_clk               ),
  .S03_AXI_araddr           (dsa_0_m_axi_araddr      ),
  .S03_AXI_arburst          (dsa_0_m_axi_arburst     ),
  .S03_AXI_arcache          (dsa_0_m_axi_arcache     ),
  .S03_AXI_aresetn          (dsa_0_rstn              ),
  .S03_AXI_arid             (dsa_0_m_axi_arid        ),
  .S03_AXI_arlen            (dsa_0_m_axi_arlen       ),
  .S03_AXI_arlock           (dsa_0_m_axi_arlock      ),
  .S03_AXI_arprot           (dsa_0_m_axi_arprot      ),
  .S03_AXI_arqos            (dsa_0_m_axi_arqos       ),
  .S03_AXI_arready          (dsa_0_m_axi_arready     ),
  .S03_AXI_arsize           (dsa_0_m_axi_arsize      ),
  .S03_AXI_arvalid          (dsa_0_m_axi_arvalid     ),
  .S03_AXI_awaddr           (dsa_0_m_axi_awaddr      ),
  .S03_AXI_awburst          (dsa_0_m_axi_awburst     ),
  .S03_AXI_awcache          (dsa_0_m_axi_awcache     ),
  .S03_AXI_awid             (dsa_0_m_axi_awid        ),
  .S03_AXI_awlen            (dsa_0_m_axi_awlen       ),
  .S03_AXI_awlock           (dsa_0_m_axi_awlock      ),
  .S03_AXI_awprot           (dsa_0_m_axi_awprot      ),
  .S03_AXI_awqos            (dsa_0_m_axi_awqos       ),
  .S03_AXI_awready          (dsa_0_m_axi_awready     ),
  .S03_AXI_awsize           (dsa_0_m_axi_awsize      ),
  .S03_AXI_awvalid          (dsa_0_m_axi_awvalid     ),
  .S03_AXI_bid              (dsa_0_m_axi_bid         ),
  .S03_AXI_bready           (dsa_0_m_axi_bready      ),
  .S03_AXI_bresp            (dsa_0_m_axi_bresp       ),
  .S03_AXI_bvalid           (dsa_0_m_axi_bvalid      ),
  .S03_AXI_rdata            (dsa_0_m_axi_rdata       ),
  .S03_AXI_rid              (dsa_0_m_axi_rid         ),
  .S03_AXI_rlast            (dsa_0_m_axi_rlast       ),
  .S03_AXI_rready           (dsa_0_m_axi_rready      ),
  .S03_AXI_rresp            (dsa_0_m_axi_rresp       ),
  .S03_AXI_rvalid           (dsa_0_m_axi_rvalid      ),
  .S03_AXI_wdata            (dsa_0_m_axi_wdata       ),
  .S03_AXI_wlast            (dsa_0_m_axi_wlast       ),
  .S03_AXI_wready           (dsa_0_m_axi_wready      ),
  .S03_AXI_wstrb            (dsa_0_m_axi_wstrb       ),
  .S03_AXI_wvalid           (dsa_0_m_axi_wvalid      ),
  .S04_AXI_aclk             (dsa_1_clk               ),
  .S04_AXI_araddr           (dsa_1_m_axi_araddr      ),
  .S04_AXI_arburst          (dsa_1_m_axi_arburst     ),
  .S04_AXI_arcache          (dsa_1_m_axi_arcache     ),
  .S04_AXI_aresetn          (dsa_1_rstn              ),
  .S04_AXI_arid             (dsa_1_m_axi_arid        ),
  .S04_AXI_arlen            (dsa_1_m_axi_arlen       ),
  .S04_AXI_arlock           (dsa_1_m_axi_arlock      ),
  .S04_AXI_arprot           (dsa_1_m_axi_arprot      ),
  .S04_AXI_arqos            (dsa_1_m_axi_arqos       ),
  .S04_AXI_arready          (dsa_1_m_axi_arready     ),
  .S04_AXI_arsize           (dsa_1_m_axi_arsize      ),
  .S04_AXI_arvalid          (dsa_1_m_axi_arvalid     ),
  .S04_AXI_awaddr           (dsa_1_m_axi_awaddr      ),
  .S04_AXI_awburst          (dsa_1_m_axi_awburst     ),
  .S04_AXI_awcache          (dsa_1_m_axi_awcache     ),
  .S04_AXI_awid             (dsa_1_m_axi_awid        ),
  .S04_AXI_awlen            (dsa_1_m_axi_awlen       ),
  .S04_AXI_awlock           (dsa_1_m_axi_awlock      ),
  .S04_AXI_awprot           (dsa_1_m_axi_awprot      ),
  .S04_AXI_awqos            (dsa_1_m_axi_awqos       ),
  .S04_AXI_awready          (dsa_1_m_axi_awready     ),
  .S04_AXI_awsize           (dsa_1_m_axi_awsize      ),
  .S04_AXI_awvalid          (dsa_1_m_axi_awvalid     ),
  .S04_AXI_bid              (dsa_1_m_axi_bid         ),
  .S04_AXI_bready           (dsa_1_m_axi_bready      ),
  .S04_AXI_bresp            (dsa_1_m_axi_bresp       ),
  .S04_AXI_bvalid           (dsa_1_m_axi_bvalid      ),
  .S04_AXI_rdata            (dsa_1_m_axi_rdata       ),
  .S04_AXI_rid              (dsa_1_m_axi_rid         ),
  .S04_AXI_rlast            (dsa_1_m_axi_rlast       ),
  .S04_AXI_rready           (dsa_1_m_axi_rready      ),
  .S04_AXI_rresp            (dsa_1_m_axi_rresp       ),
  .S04_AXI_rvalid           (dsa_1_m_axi_rvalid      ),
  .S04_AXI_wdata            (dsa_1_m_axi_wdata       ),
  .S04_AXI_wlast            (dsa_1_m_axi_wlast       ),
  .S04_AXI_wready           (dsa_1_m_axi_wready      ),
  .S04_AXI_wstrb            (dsa_1_m_axi_wstrb       ),
  .S04_AXI_wvalid           (dsa_1_m_axi_wvalid      ),
  .S05_AXI_aclk             (dsa_2_clk               ),
  .S05_AXI_araddr           (dsa_2_m_axi_araddr      ),
  .S05_AXI_arburst          (dsa_2_m_axi_arburst     ),
  .S05_AXI_arcache          (dsa_2_m_axi_arcache     ),
  .S05_AXI_aresetn          (dsa_2_rstn              ),
  .S05_AXI_arid             (dsa_2_m_axi_arid        ),
  .S05_AXI_arlen            (dsa_2_m_axi_arlen       ),
  .S05_AXI_arlock           (dsa_2_m_axi_arlock      ),
  .S05_AXI_arprot           (dsa_2_m_axi_arprot      ),
  .S05_AXI_arqos            (dsa_2_m_axi_arqos       ),
  .S05_AXI_arready          (dsa_2_m_axi_arready     ),
  .S05_AXI_arsize           (dsa_2_m_axi_arsize      ),
  .S05_AXI_arvalid          (dsa_2_m_axi_arvalid     ),
  .S05_AXI_awaddr           (dsa_2_m_axi_awaddr      ),
  .S05_AXI_awburst          (dsa_2_m_axi_awburst     ),
  .S05_AXI_awcache          (dsa_2_m_axi_awcache     ),
  .S05_AXI_awid             (dsa_2_m_axi_awid        ),
  .S05_AXI_awlen            (dsa_2_m_axi_awlen       ),
  .S05_AXI_awlock           (dsa_2_m_axi_awlock      ),
  .S05_AXI_awprot           (dsa_2_m_axi_awprot      ),
  .S05_AXI_awqos            (dsa_2_m_axi_awqos       ),
  .S05_AXI_awready          (dsa_2_m_axi_awready     ),
  .S05_AXI_awsize           (dsa_2_m_axi_awsize      ),
  .S05_AXI_awvalid          (dsa_2_m_axi_awvalid     ),
  .S05_AXI_bid              (dsa_2_m_axi_bid         ),
  .S05_AXI_bready           (dsa_2_m_axi_bready      ),
  .S05_AXI_bresp            (dsa_2_m_axi_bresp       ),
  .S05_AXI_bvalid           (dsa_2_m_axi_bvalid      ),
  .S05_AXI_rdata            (dsa_2_m_axi_rdata       ),
  .S05_AXI_rid              (dsa_2_m_axi_rid         ),
  .S05_AXI_rlast            (dsa_2_m_axi_rlast       ),
  .S05_AXI_rready           (dsa_2_m_axi_rready      ),
  .S05_AXI_rresp            (dsa_2_m_axi_rresp       ),
  .S05_AXI_rvalid           (dsa_2_m_axi_rvalid      ),
  .S05_AXI_wdata            (dsa_2_m_axi_wdata       ),
  .S05_AXI_wlast            (dsa_2_m_axi_wlast       ),
  .S05_AXI_wready           (dsa_2_m_axi_wready      ),
  .S05_AXI_wstrb            (dsa_2_m_axi_wstrb       ),
  .S05_AXI_wvalid           (dsa_2_m_axi_wvalid      )
);

// &Connect( @65
//     .S00_AXI_aclk (rv_0_clk), @66
//     .S00_AXI_aresetn (rv_0_rstn), @67
//     .S01_AXI_aclk (rv_1_clk), @68
//     .S01_AXI_aresetn (rv_1_rstn), @69
//     .S02_AXI_aclk (rv_2_clk), @70
//     .S02_AXI_aresetn (rv_2_rstn), @71
//     .S03_AXI_aclk (dsa_0_clk), @72
//     .S03_AXI_aresetn (dsa_0_rstn), @73
//     .S04_AXI_aclk (dsa_1_clk), @74
//     .S04_AXI_aresetn (dsa_1_rstn), @75
//     .S05_AXI_aclk (dsa_2_clk), @76
//     .S05_AXI_aresetn (dsa_2_rstn), @77
//     .M00_AXI_aclk (mem_sub_sys_clk), @78
//     .M00_AXI_aresetn (mem_sub_sys_rstn), @79
//     .M01_AXI_aclk (mem_sub_sys_clk), @80
//     .M01_AXI_aresetn (mem_sub_sys_rstn), @81
//     .M02_AXI_aclk (mem_sub_sys_clk), @82
//     .M02_AXI_aresetn (mem_sub_sys_rstn), @83
//     .M03_AXI_aclk (mem_sub_sys_clk), @84
//     .M03_AXI_aresetn (mem_sub_sys_rstn), @85
// ); @86

// &ModuleEnd; @88
endmodule


