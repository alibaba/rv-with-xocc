/* 
*Copyright (c) 2021, Alibaba Group;
*Licensed under the Apache License, Version 2.0 (the "License");
*you may not use this file except in compliance with the License.
*You may obtain a copy of the License at

*   http://www.apache.org/licenses/LICENSE-2.0

*Unless required by applicable law or agreed to in writing, software
*distributed under the License is distributed on an "AS IS" BASIS,
*WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
*See the License for the specific language governing permissions and
*limitations under the License.
*/

// SPM Memory Initialization  
defparam `PE_0_0_SPM.x_axi_uram_0.MEMORY_INIT_FILE="pe_0_0_mem_0_init.mem";
defparam `PE_0_0_SPM.x_axi_uram_1.MEMORY_INIT_FILE="pe_0_0_mem_1_init.mem";
defparam `PE_0_0_SPM.x_axi_uram_2.MEMORY_INIT_FILE="pe_0_0_mem_2_init.mem";
defparam `PE_0_0_SPM.x_axi_uram_3.MEMORY_INIT_FILE="pe_0_0_mem_3_init.mem";

